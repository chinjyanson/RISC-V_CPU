module ALU_top #(
    parameter DATA_WIDTH = 32 
)(
    input 
)