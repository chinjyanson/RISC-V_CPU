module maindecoder #(
    parameters  OP_WIDTH = 7,
    parameters  IMM_WIDTH = 2
) (
    port_list
);
    
endmodule