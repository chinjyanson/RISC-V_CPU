heye heye




