module aludecoder #(


)(
    input   logic [OP_WIDTH-1:0]    opcode_i,
    output  logic []
);
    
endmodule