module top (
    input logic         clk,
    input logic         rst,
    output logic        anot0
);






