module controller #(
    parameters OP_WIDTH = 7
) (
    input   logic                   clk,
    input   logic [OP_WIDTH-1:0]    op,
    input   logic
);
    
endmodule