/*
	Function: Control Unit Pipeline Register between Instruction Execution and Memory Access Stage
*/