module alu (
    input logic [2:0] ALUControl,
    input logic [31:0] SrcA,
    input logic [31:0] SrcB,
    
)