module name #(
    parameters  OP_WIDTH = 7,
    parameters  IMM_WIDTH = 2

)(
    input   logic [OP_WIDTH-1:0]    opcode_i,
    output  logic []
);
    
endmodule