module red_top #(
    parameter DATA_WIDTH = 32 
)(
    input wire 
)

endmodule
