module controller #(
    parameters
) (
    port_list
);
    
endmodule